NAND2 cell simulation
.include "./lib/prelude.spice"

* include target cell model
.include "./sky130_fd_sc_hd/cells/nand2/sky130_fd_sc_hd__nand2_8.spice"

* create target cell
xcell A B Vgnd Vgnd Vdd Vdd Y sky130_fd_sc_hd__nand2_8

* set gnd and power
Vgnd Vgnd 0 0
Vdd Vdd Vgnd 1.8

* create test pulses
Va A Vgnd pulse(0 1.8 1n 10p 10p 1n 2n)
Vb B Vgnd pulse(0 1.8 1.5n 10p 10p 1n 2n)

* setup the transient analysis
.tran 10p 3n 0

.control
run

hardcopy plots/nand_2.ps A B Y
shell open plots/nand_2.ps

exit
.endc