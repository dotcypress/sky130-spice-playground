.lib "./sky130_fd_pr/models/sky130.lib.spice" tt

.control
set hcopydevtype=postscript
set hcopypscolor=1
set hcopywidth=1280
set hcopyheight=720
.endc

.end
